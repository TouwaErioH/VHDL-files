library verilog;
use verilog.vl_types.all;
entity pipecomp_tb is
end pipecomp_tb;
