library verilog;
use verilog.vl_types.all;
entity plcomp_tb is
end plcomp_tb;
